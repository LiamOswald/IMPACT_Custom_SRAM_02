VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO full_sram
  CLASS BLOCK ;
  FOREIGN full_sram ;
  ORIGIN 23.200 1875.000 ;
  SIZE 251.200 BY 1908.000 ;
  PIN DataIn0
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 1.250 -1875.000 2.200 -1873.000 ;
    END
  END DataIn0
  PIN DataOut0
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 4.800 -1875.000 5.400 -1873.000 ;
    END
  END DataOut0
  PIN DataIn1
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 8.050 -1875.000 9.000 -1873.000 ;
    END
  END DataIn1
  PIN DataOut1
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 11.650 -1875.000 12.250 -1873.000 ;
    END
  END DataOut1
  PIN DataIn2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 14.850 -1875.000 15.800 -1873.000 ;
    END
  END DataIn2
  PIN DataOut2
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 18.400 -1875.000 19.000 -1873.000 ;
    END
  END DataOut2
  PIN DataIn3
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 21.650 -1875.000 22.600 -1873.000 ;
    END
  END DataIn3
  PIN DataOut3
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 25.150 -1875.000 25.750 -1873.000 ;
    END
  END DataOut3
  PIN DataIn4
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 28.450 -1875.000 29.400 -1873.000 ;
    END
  END DataIn4
  PIN DataOut4
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 31.900 -1875.000 32.500 -1873.000 ;
    END
  END DataOut4
  PIN DataIn5
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 35.250 -1875.000 36.200 -1873.000 ;
    END
  END DataIn5
  PIN DataOut5
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 38.650 -1875.000 39.250 -1873.000 ;
    END
  END DataOut5
  PIN DataIn6
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 42.050 -1875.000 43.000 -1873.000 ;
    END
  END DataIn6
  PIN DataOut6
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 45.400 -1875.000 46.000 -1873.000 ;
    END
  END DataOut6
  PIN DataIn7
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 -1875.000 49.800 -1873.000 ;
    END
  END DataIn7
  PIN DataOut7
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 52.150 -1875.000 52.750 -1873.000 ;
    END
  END DataOut7
  PIN DataIn8
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 55.650 -1875.000 56.600 -1873.000 ;
    END
  END DataIn8
  PIN DataOut8
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 58.900 -1875.000 59.500 -1873.000 ;
    END
  END DataOut8
  PIN DataIn9
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 62.450 -1875.000 63.400 -1873.000 ;
    END
  END DataIn9
  PIN DataOut9
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 65.650 -1875.000 66.250 -1873.000 ;
    END
  END DataOut9
  PIN DataIn10
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 69.250 -1875.000 70.200 -1873.000 ;
    END
  END DataIn10
  PIN DataOut10
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 72.400 -1875.000 73.000 -1873.000 ;
    END
  END DataOut10
  PIN DataIn11
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 76.050 -1875.000 77.000 -1873.000 ;
    END
  END DataIn11
  PIN DataOut11
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 79.150 -1875.000 79.750 -1873.000 ;
    END
  END DataOut11
  PIN DataIn12
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 82.850 -1875.000 83.800 -1873.000 ;
    END
  END DataIn12
  PIN DataOut12
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 85.900 -1875.000 86.500 -1873.000 ;
    END
  END DataOut12
  PIN DataIn13
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 89.650 -1875.000 90.600 -1873.000 ;
    END
  END DataIn13
  PIN DataOut13
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 92.650 -1875.000 93.250 -1873.000 ;
    END
  END DataOut13
  PIN DataIn14
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 96.450 -1875.000 97.400 -1873.000 ;
    END
  END DataIn14
  PIN DataOut14
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 99.400 -1875.000 100.000 -1873.000 ;
    END
  END DataOut14
  PIN DataIn15
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 103.250 -1875.000 104.200 -1873.000 ;
    END
  END DataIn15
  PIN DataOut15
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 106.150 -1875.000 106.750 -1873.000 ;
    END
  END DataOut15
  PIN DataIn16
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 110.050 -1875.000 111.000 -1873.000 ;
    END
  END DataIn16
  PIN DataOut16
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 112.900 -1875.000 113.500 -1873.000 ;
    END
  END DataOut16
  PIN DataIn17
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 116.850 -1875.000 117.800 -1873.000 ;
    END
  END DataIn17
  PIN DataOut17
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 119.650 -1875.000 120.250 -1873.000 ;
    END
  END DataOut17
  PIN DataIn18
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 123.650 -1875.000 124.600 -1873.000 ;
    END
  END DataIn18
  PIN DataOut18
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 126.400 -1875.000 127.000 -1873.000 ;
    END
  END DataOut18
  PIN DataIn19
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 130.450 -1875.000 131.400 -1873.000 ;
    END
  END DataIn19
  PIN DataOut19
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 133.150 -1875.000 133.750 -1873.000 ;
    END
  END DataOut19
  PIN DataIn20
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 137.250 -1875.000 138.200 -1873.000 ;
    END
  END DataIn20
  PIN DataOut20
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 139.900 -1875.000 140.500 -1873.000 ;
    END
  END DataOut20
  PIN DataIn21
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 144.050 -1875.000 145.000 -1873.000 ;
    END
  END DataIn21
  PIN DataOut21
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 146.650 -1875.000 147.250 -1873.000 ;
    END
  END DataOut21
  PIN DataIn22
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 150.850 -1875.000 151.800 -1873.000 ;
    END
  END DataIn22
  PIN DataOut22
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 153.400 -1875.000 154.000 -1873.000 ;
    END
  END DataOut22
  PIN DataIn23
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 157.650 -1875.000 158.600 -1873.000 ;
    END
  END DataIn23
  PIN DataOut23
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 160.150 -1875.000 160.750 -1873.000 ;
    END
  END DataOut23
  PIN DataIn24
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 164.450 -1875.000 165.400 -1873.000 ;
    END
  END DataIn24
  PIN DataOut24
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 166.900 -1875.000 167.500 -1873.000 ;
    END
  END DataOut24
  PIN DataIn25
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 171.250 -1875.000 172.200 -1873.000 ;
    END
  END DataIn25
  PIN DataOut25
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 173.650 -1875.000 174.250 -1873.000 ;
    END
  END DataOut25
  PIN DataIn26
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 178.050 -1875.000 179.000 -1873.000 ;
    END
  END DataIn26
  PIN DataOut26
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 180.400 -1875.000 181.000 -1873.000 ;
    END
  END DataOut26
  PIN DataIn27
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 184.850 -1875.000 185.800 -1873.000 ;
    END
  END DataIn27
  PIN DataOut27
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 187.150 -1875.000 187.750 -1873.000 ;
    END
  END DataOut27
  PIN DataIn28
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 191.650 -1875.000 192.600 -1873.000 ;
    END
  END DataIn28
  PIN DataOut28
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 193.900 -1875.000 194.500 -1873.000 ;
    END
  END DataOut28
  PIN DataIn29
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 198.450 -1875.000 199.400 -1873.000 ;
    END
  END DataIn29
  PIN DataOut29
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 200.650 -1875.000 201.250 -1873.000 ;
    END
  END DataOut29
  PIN DataIn30
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 205.250 -1875.000 206.200 -1873.000 ;
    END
  END DataIn30
  PIN DataOut30
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 207.400 -1875.000 208.000 -1873.000 ;
    END
  END DataOut30
  PIN DataIn31
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met2 ;
        RECT 212.050 -1875.000 213.000 -1873.000 ;
    END
  END DataIn31
  PIN DataOut31
    ANTENNADIFFAREA 0.411600 ;
    PORT
      LAYER met2 ;
        RECT 214.150 -1875.000 214.750 -1873.000 ;
    END
  END DataOut31
  PIN writeen
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1851.450 -21.200 -1850.450 ;
    END
  END writeen
  PIN readen
    ANTENNAGATEAREA 7.257600 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1838.950 -21.200 -1837.950 ;
    END
  END readen
  PIN PRE
    ANTENNAGATEAREA 8.294400 ;
    PORT
      LAYER met3 ;
        RECT -23.200 20.450 -21.200 21.450 ;
    END
  END PRE
  PIN WL0
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 15.250 -21.200 16.250 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 13.900 -21.200 14.900 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 11.650 -21.200 12.650 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 10.300 -21.200 11.300 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 8.050 -21.200 9.050 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 6.700 -21.200 7.700 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 4.450 -21.200 5.450 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 3.100 -21.200 4.100 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 0.850 -21.200 1.850 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -0.500 -21.200 0.500 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -2.750 -21.200 -1.750 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -4.100 -21.200 -3.100 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -6.350 -21.200 -5.350 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -7.700 -21.200 -6.700 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -9.950 -21.200 -8.950 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -11.300 -21.200 -10.300 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -13.550 -21.200 -12.550 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -14.900 -21.200 -13.900 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -17.150 -21.200 -16.150 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -18.500 -21.200 -17.500 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -20.750 -21.200 -19.750 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -22.100 -21.200 -21.100 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -24.350 -21.200 -23.350 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -25.700 -21.200 -24.700 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -27.950 -21.200 -26.950 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -29.300 -21.200 -28.300 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -31.550 -21.200 -30.550 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -32.900 -21.200 -31.900 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -35.150 -21.200 -34.150 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -36.500 -21.200 -35.500 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -38.750 -21.200 -37.750 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -40.100 -21.200 -39.100 ;
    END
  END WL31
  PIN WL32
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -42.350 -21.200 -41.350 ;
    END
  END WL32
  PIN WL33
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -43.700 -21.200 -42.700 ;
    END
  END WL33
  PIN WL34
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -45.950 -21.200 -44.950 ;
    END
  END WL34
  PIN WL35
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -47.300 -21.200 -46.300 ;
    END
  END WL35
  PIN WL36
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -49.550 -21.200 -48.550 ;
    END
  END WL36
  PIN WL37
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -50.900 -21.200 -49.900 ;
    END
  END WL37
  PIN WL38
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -53.150 -21.200 -52.150 ;
    END
  END WL38
  PIN WL39
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -54.500 -21.200 -53.500 ;
    END
  END WL39
  PIN WL40
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -56.750 -21.200 -55.750 ;
    END
  END WL40
  PIN WL41
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -58.100 -21.200 -57.100 ;
    END
  END WL41
  PIN WL42
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -60.350 -21.200 -59.350 ;
    END
  END WL42
  PIN WL43
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -61.700 -21.200 -60.700 ;
    END
  END WL43
  PIN WL44
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -63.950 -21.200 -62.950 ;
    END
  END WL44
  PIN WL45
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -65.300 -21.200 -64.300 ;
    END
  END WL45
  PIN WL46
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -67.550 -21.200 -66.550 ;
    END
  END WL46
  PIN WL47
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -68.900 -21.200 -67.900 ;
    END
  END WL47
  PIN WL48
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -71.150 -21.200 -70.150 ;
    END
  END WL48
  PIN WL49
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -72.500 -21.200 -71.500 ;
    END
  END WL49
  PIN WL50
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -74.750 -21.200 -73.750 ;
    END
  END WL50
  PIN WL51
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -76.100 -21.200 -75.100 ;
    END
  END WL51
  PIN WL52
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -78.350 -21.200 -77.350 ;
    END
  END WL52
  PIN WL53
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -79.700 -21.200 -78.700 ;
    END
  END WL53
  PIN WL54
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -81.950 -21.200 -80.950 ;
    END
  END WL54
  PIN WL55
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -83.300 -21.200 -82.300 ;
    END
  END WL55
  PIN WL56
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -85.550 -21.200 -84.550 ;
    END
  END WL56
  PIN WL57
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -86.900 -21.200 -85.900 ;
    END
  END WL57
  PIN WL58
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -89.150 -21.200 -88.150 ;
    END
  END WL58
  PIN WL59
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -90.500 -21.200 -89.500 ;
    END
  END WL59
  PIN WL60
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -92.750 -21.200 -91.750 ;
    END
  END WL60
  PIN WL61
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -94.100 -21.200 -93.100 ;
    END
  END WL61
  PIN WL62
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -96.350 -21.200 -95.350 ;
    END
  END WL62
  PIN WL63
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -97.700 -21.200 -96.700 ;
    END
  END WL63
  PIN WL64
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -99.950 -21.200 -98.950 ;
    END
  END WL64
  PIN WL65
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -101.300 -21.200 -100.300 ;
    END
  END WL65
  PIN WL66
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -103.550 -21.200 -102.550 ;
    END
  END WL66
  PIN WL67
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -104.900 -21.200 -103.900 ;
    END
  END WL67
  PIN WL68
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -107.150 -21.200 -106.150 ;
    END
  END WL68
  PIN WL69
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -108.500 -21.200 -107.500 ;
    END
  END WL69
  PIN WL70
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -110.750 -21.200 -109.750 ;
    END
  END WL70
  PIN WL71
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -112.100 -21.200 -111.100 ;
    END
  END WL71
  PIN WL72
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -114.350 -21.200 -113.350 ;
    END
  END WL72
  PIN WL73
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -115.700 -21.200 -114.700 ;
    END
  END WL73
  PIN WL74
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -117.950 -21.200 -116.950 ;
    END
  END WL74
  PIN WL75
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -119.300 -21.200 -118.300 ;
    END
  END WL75
  PIN WL76
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -121.550 -21.200 -120.550 ;
    END
  END WL76
  PIN WL77
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -122.900 -21.200 -121.900 ;
    END
  END WL77
  PIN WL78
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -125.150 -21.200 -124.150 ;
    END
  END WL78
  PIN WL79
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -126.500 -21.200 -125.500 ;
    END
  END WL79
  PIN WL80
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -128.750 -21.200 -127.750 ;
    END
  END WL80
  PIN WL81
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -130.100 -21.200 -129.100 ;
    END
  END WL81
  PIN WL82
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -132.350 -21.200 -131.350 ;
    END
  END WL82
  PIN WL83
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -133.700 -21.200 -132.700 ;
    END
  END WL83
  PIN WL84
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -135.950 -21.200 -134.950 ;
    END
  END WL84
  PIN WL85
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -137.300 -21.200 -136.300 ;
    END
  END WL85
  PIN WL86
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -139.550 -21.200 -138.550 ;
    END
  END WL86
  PIN WL87
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -140.900 -21.200 -139.900 ;
    END
  END WL87
  PIN WL88
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -143.150 -21.200 -142.150 ;
    END
  END WL88
  PIN WL89
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -144.500 -21.200 -143.500 ;
    END
  END WL89
  PIN WL90
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -146.750 -21.200 -145.750 ;
    END
  END WL90
  PIN WL91
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -148.100 -21.200 -147.100 ;
    END
  END WL91
  PIN WL92
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -150.350 -21.200 -149.350 ;
    END
  END WL92
  PIN WL93
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -151.700 -21.200 -150.700 ;
    END
  END WL93
  PIN WL94
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -153.950 -21.200 -152.950 ;
    END
  END WL94
  PIN WL95
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -155.300 -21.200 -154.300 ;
    END
  END WL95
  PIN WL96
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -157.550 -21.200 -156.550 ;
    END
  END WL96
  PIN WL97
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -158.900 -21.200 -157.900 ;
    END
  END WL97
  PIN WL98
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -161.150 -21.200 -160.150 ;
    END
  END WL98
  PIN WL99
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -162.500 -21.200 -161.500 ;
    END
  END WL99
  PIN WL100
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -164.750 -21.200 -163.750 ;
    END
  END WL100
  PIN WL101
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -166.100 -21.200 -165.100 ;
    END
  END WL101
  PIN WL102
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -168.350 -21.200 -167.350 ;
    END
  END WL102
  PIN WL103
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -169.700 -21.200 -168.700 ;
    END
  END WL103
  PIN WL104
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -171.950 -21.200 -170.950 ;
    END
  END WL104
  PIN WL105
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -173.300 -21.200 -172.300 ;
    END
  END WL105
  PIN WL106
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -175.550 -21.200 -174.550 ;
    END
  END WL106
  PIN WL107
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -176.900 -21.200 -175.900 ;
    END
  END WL107
  PIN WL108
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -179.150 -21.200 -178.150 ;
    END
  END WL108
  PIN WL109
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -180.500 -21.200 -179.500 ;
    END
  END WL109
  PIN WL110
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -182.750 -21.200 -181.750 ;
    END
  END WL110
  PIN WL111
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -184.100 -21.200 -183.100 ;
    END
  END WL111
  PIN WL112
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -186.350 -21.200 -185.350 ;
    END
  END WL112
  PIN WL113
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -187.700 -21.200 -186.700 ;
    END
  END WL113
  PIN WL114
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -190.500 -21.200 -189.500 ;
    END
  END WL114
  PIN WL115
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -191.850 -21.200 -190.850 ;
    END
  END WL115
  PIN WL116
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -194.100 -21.200 -193.100 ;
    END
  END WL116
  PIN WL117
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -195.450 -21.200 -194.450 ;
    END
  END WL117
  PIN WL118
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -197.700 -21.200 -196.700 ;
    END
  END WL118
  PIN WL119
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -199.050 -21.200 -198.050 ;
    END
  END WL119
  PIN WL120
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -201.300 -21.200 -200.300 ;
    END
  END WL120
  PIN WL121
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -202.650 -21.200 -201.650 ;
    END
  END WL121
  PIN WL122
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -204.900 -21.200 -203.900 ;
    END
  END WL122
  PIN WL123
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -206.250 -21.200 -205.250 ;
    END
  END WL123
  PIN WL124
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -208.500 -21.200 -207.500 ;
    END
  END WL124
  PIN WL125
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -209.850 -21.200 -208.850 ;
    END
  END WL125
  PIN WL126
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -212.100 -21.200 -211.100 ;
    END
  END WL126
  PIN WL127
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -213.450 -21.200 -212.450 ;
    END
  END WL127
  PIN WL128
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -215.700 -21.200 -214.700 ;
    END
  END WL128
  PIN WL129
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -217.050 -21.200 -216.050 ;
    END
  END WL129
  PIN WL130
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -219.300 -21.200 -218.300 ;
    END
  END WL130
  PIN WL131
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -220.650 -21.200 -219.650 ;
    END
  END WL131
  PIN WL132
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -222.900 -21.200 -221.900 ;
    END
  END WL132
  PIN WL133
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -224.250 -21.200 -223.250 ;
    END
  END WL133
  PIN WL134
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -226.500 -21.200 -225.500 ;
    END
  END WL134
  PIN WL135
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -227.850 -21.200 -226.850 ;
    END
  END WL135
  PIN WL136
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -230.100 -21.200 -229.100 ;
    END
  END WL136
  PIN WL137
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -231.450 -21.200 -230.450 ;
    END
  END WL137
  PIN WL138
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -233.700 -21.200 -232.700 ;
    END
  END WL138
  PIN WL139
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -235.050 -21.200 -234.050 ;
    END
  END WL139
  PIN WL140
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -237.300 -21.200 -236.300 ;
    END
  END WL140
  PIN WL141
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -238.650 -21.200 -237.650 ;
    END
  END WL141
  PIN WL142
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -240.900 -21.200 -239.900 ;
    END
  END WL142
  PIN WL143
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -242.250 -21.200 -241.250 ;
    END
  END WL143
  PIN WL144
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -244.500 -21.200 -243.500 ;
    END
  END WL144
  PIN WL145
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -245.850 -21.200 -244.850 ;
    END
  END WL145
  PIN WL146
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -248.100 -21.200 -247.100 ;
    END
  END WL146
  PIN WL147
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -249.450 -21.200 -248.450 ;
    END
  END WL147
  PIN WL148
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -251.700 -21.200 -250.700 ;
    END
  END WL148
  PIN WL149
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -253.050 -21.200 -252.050 ;
    END
  END WL149
  PIN WL150
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -255.300 -21.200 -254.300 ;
    END
  END WL150
  PIN WL151
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -256.650 -21.200 -255.650 ;
    END
  END WL151
  PIN WL152
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -258.900 -21.200 -257.900 ;
    END
  END WL152
  PIN WL153
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -260.250 -21.200 -259.250 ;
    END
  END WL153
  PIN WL154
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -262.500 -21.200 -261.500 ;
    END
  END WL154
  PIN WL155
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -263.850 -21.200 -262.850 ;
    END
  END WL155
  PIN WL156
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -266.100 -21.200 -265.100 ;
    END
  END WL156
  PIN WL157
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -267.450 -21.200 -266.450 ;
    END
  END WL157
  PIN WL158
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -269.700 -21.200 -268.700 ;
    END
  END WL158
  PIN WL159
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -271.050 -21.200 -270.050 ;
    END
  END WL159
  PIN WL160
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -273.300 -21.200 -272.300 ;
    END
  END WL160
  PIN WL161
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -274.650 -21.200 -273.650 ;
    END
  END WL161
  PIN WL162
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -276.900 -21.200 -275.900 ;
    END
  END WL162
  PIN WL163
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -278.250 -21.200 -277.250 ;
    END
  END WL163
  PIN WL164
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -280.500 -21.200 -279.500 ;
    END
  END WL164
  PIN WL165
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -281.850 -21.200 -280.850 ;
    END
  END WL165
  PIN WL166
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -284.100 -21.200 -283.100 ;
    END
  END WL166
  PIN WL167
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -285.450 -21.200 -284.450 ;
    END
  END WL167
  PIN WL168
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -287.700 -21.200 -286.700 ;
    END
  END WL168
  PIN WL169
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -289.050 -21.200 -288.050 ;
    END
  END WL169
  PIN WL170
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -291.300 -21.200 -290.300 ;
    END
  END WL170
  PIN WL171
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -292.650 -21.200 -291.650 ;
    END
  END WL171
  PIN WL172
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -294.900 -21.200 -293.900 ;
    END
  END WL172
  PIN WL173
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -296.250 -21.200 -295.250 ;
    END
  END WL173
  PIN WL174
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -298.500 -21.200 -297.500 ;
    END
  END WL174
  PIN WL175
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -299.850 -21.200 -298.850 ;
    END
  END WL175
  PIN WL176
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -302.100 -21.200 -301.100 ;
    END
  END WL176
  PIN WL177
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -303.450 -21.200 -302.450 ;
    END
  END WL177
  PIN WL178
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -305.700 -21.200 -304.700 ;
    END
  END WL178
  PIN WL179
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -307.050 -21.200 -306.050 ;
    END
  END WL179
  PIN WL180
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -309.300 -21.200 -308.300 ;
    END
  END WL180
  PIN WL181
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -310.650 -21.200 -309.650 ;
    END
  END WL181
  PIN WL182
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -312.900 -21.200 -311.900 ;
    END
  END WL182
  PIN WL183
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -314.250 -21.200 -313.250 ;
    END
  END WL183
  PIN WL184
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -316.500 -21.200 -315.500 ;
    END
  END WL184
  PIN WL185
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -317.850 -21.200 -316.850 ;
    END
  END WL185
  PIN WL186
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -320.100 -21.200 -319.100 ;
    END
  END WL186
  PIN WL187
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -321.450 -21.200 -320.450 ;
    END
  END WL187
  PIN WL188
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -323.700 -21.200 -322.700 ;
    END
  END WL188
  PIN WL189
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -325.050 -21.200 -324.050 ;
    END
  END WL189
  PIN WL190
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -327.300 -21.200 -326.300 ;
    END
  END WL190
  PIN WL191
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -328.650 -21.200 -327.650 ;
    END
  END WL191
  PIN WL192
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -330.900 -21.200 -329.900 ;
    END
  END WL192
  PIN WL193
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -332.250 -21.200 -331.250 ;
    END
  END WL193
  PIN WL194
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -334.500 -21.200 -333.500 ;
    END
  END WL194
  PIN WL195
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -335.850 -21.200 -334.850 ;
    END
  END WL195
  PIN WL196
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -338.100 -21.200 -337.100 ;
    END
  END WL196
  PIN WL197
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -339.450 -21.200 -338.450 ;
    END
  END WL197
  PIN WL198
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -341.700 -21.200 -340.700 ;
    END
  END WL198
  PIN WL199
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -343.050 -21.200 -342.050 ;
    END
  END WL199
  PIN WL200
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -345.300 -21.200 -344.300 ;
    END
  END WL200
  PIN WL201
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -346.650 -21.200 -345.650 ;
    END
  END WL201
  PIN WL202
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -348.900 -21.200 -347.900 ;
    END
  END WL202
  PIN WL203
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -350.250 -21.200 -349.250 ;
    END
  END WL203
  PIN WL204
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -352.500 -21.200 -351.500 ;
    END
  END WL204
  PIN WL205
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -353.850 -21.200 -352.850 ;
    END
  END WL205
  PIN WL206
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -356.100 -21.200 -355.100 ;
    END
  END WL206
  PIN WL207
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -357.450 -21.200 -356.450 ;
    END
  END WL207
  PIN WL208
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -359.700 -21.200 -358.700 ;
    END
  END WL208
  PIN WL209
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -361.050 -21.200 -360.050 ;
    END
  END WL209
  PIN WL210
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -363.300 -21.200 -362.300 ;
    END
  END WL210
  PIN WL211
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -364.650 -21.200 -363.650 ;
    END
  END WL211
  PIN WL212
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -366.900 -21.200 -365.900 ;
    END
  END WL212
  PIN WL213
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -368.250 -21.200 -367.250 ;
    END
  END WL213
  PIN WL214
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -370.500 -21.200 -369.500 ;
    END
  END WL214
  PIN WL215
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -371.850 -21.200 -370.850 ;
    END
  END WL215
  PIN WL216
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -374.100 -21.200 -373.100 ;
    END
  END WL216
  PIN WL217
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -375.450 -21.200 -374.450 ;
    END
  END WL217
  PIN WL218
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -377.700 -21.200 -376.700 ;
    END
  END WL218
  PIN WL219
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -379.050 -21.200 -378.050 ;
    END
  END WL219
  PIN WL220
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -381.300 -21.200 -380.300 ;
    END
  END WL220
  PIN WL221
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -382.650 -21.200 -381.650 ;
    END
  END WL221
  PIN WL222
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -384.900 -21.200 -383.900 ;
    END
  END WL222
  PIN WL223
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -386.250 -21.200 -385.250 ;
    END
  END WL223
  PIN WL224
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -389.050 -21.200 -388.050 ;
    END
  END WL224
  PIN WL225
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -390.400 -21.200 -389.400 ;
    END
  END WL225
  PIN WL226
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -392.650 -21.200 -391.650 ;
    END
  END WL226
  PIN WL227
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -394.000 -21.200 -393.000 ;
    END
  END WL227
  PIN WL228
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -396.250 -21.200 -395.250 ;
    END
  END WL228
  PIN WL229
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -397.600 -21.200 -396.600 ;
    END
  END WL229
  PIN WL230
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -399.850 -21.200 -398.850 ;
    END
  END WL230
  PIN WL231
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -401.200 -21.200 -400.200 ;
    END
  END WL231
  PIN WL232
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -403.450 -21.200 -402.450 ;
    END
  END WL232
  PIN WL233
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -404.800 -21.200 -403.800 ;
    END
  END WL233
  PIN WL234
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -407.050 -21.200 -406.050 ;
    END
  END WL234
  PIN WL235
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -408.400 -21.200 -407.400 ;
    END
  END WL235
  PIN WL236
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -410.650 -21.200 -409.650 ;
    END
  END WL236
  PIN WL237
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -412.000 -21.200 -411.000 ;
    END
  END WL237
  PIN WL238
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -414.250 -21.200 -413.250 ;
    END
  END WL238
  PIN WL239
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -415.600 -21.200 -414.600 ;
    END
  END WL239
  PIN WL240
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -417.850 -21.200 -416.850 ;
    END
  END WL240
  PIN WL241
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -419.200 -21.200 -418.200 ;
    END
  END WL241
  PIN WL242
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -421.450 -21.200 -420.450 ;
    END
  END WL242
  PIN WL243
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -422.800 -21.200 -421.800 ;
    END
  END WL243
  PIN WL244
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -425.050 -21.200 -424.050 ;
    END
  END WL244
  PIN WL245
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -426.400 -21.200 -425.400 ;
    END
  END WL245
  PIN WL246
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -428.650 -21.200 -427.650 ;
    END
  END WL246
  PIN WL247
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -430.000 -21.200 -429.000 ;
    END
  END WL247
  PIN WL248
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -432.250 -21.200 -431.250 ;
    END
  END WL248
  PIN WL249
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -433.600 -21.200 -432.600 ;
    END
  END WL249
  PIN WL250
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -435.850 -21.200 -434.850 ;
    END
  END WL250
  PIN WL251
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -437.200 -21.200 -436.200 ;
    END
  END WL251
  PIN WL252
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -439.450 -21.200 -438.450 ;
    END
  END WL252
  PIN WL253
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -440.800 -21.200 -439.800 ;
    END
  END WL253
  PIN WL254
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -443.050 -21.200 -442.050 ;
    END
  END WL254
  PIN WL255
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -444.400 -21.200 -443.400 ;
    END
  END WL255
  PIN WL256
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -446.650 -21.200 -445.650 ;
    END
  END WL256
  PIN WL257
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -448.000 -21.200 -447.000 ;
    END
  END WL257
  PIN WL258
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -450.250 -21.200 -449.250 ;
    END
  END WL258
  PIN WL259
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -451.600 -21.200 -450.600 ;
    END
  END WL259
  PIN WL260
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -453.850 -21.200 -452.850 ;
    END
  END WL260
  PIN WL261
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -455.200 -21.200 -454.200 ;
    END
  END WL261
  PIN WL262
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -457.450 -21.200 -456.450 ;
    END
  END WL262
  PIN WL263
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -458.800 -21.200 -457.800 ;
    END
  END WL263
  PIN WL264
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -461.050 -21.200 -460.050 ;
    END
  END WL264
  PIN WL265
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -462.400 -21.200 -461.400 ;
    END
  END WL265
  PIN WL266
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -464.650 -21.200 -463.650 ;
    END
  END WL266
  PIN WL267
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -466.000 -21.200 -465.000 ;
    END
  END WL267
  PIN WL268
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -468.250 -21.200 -467.250 ;
    END
  END WL268
  PIN WL269
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -469.600 -21.200 -468.600 ;
    END
  END WL269
  PIN WL270
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -471.850 -21.200 -470.850 ;
    END
  END WL270
  PIN WL271
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -473.200 -21.200 -472.200 ;
    END
  END WL271
  PIN WL272
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -475.450 -21.200 -474.450 ;
    END
  END WL272
  PIN WL273
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -476.800 -21.200 -475.800 ;
    END
  END WL273
  PIN WL274
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -479.050 -21.200 -478.050 ;
    END
  END WL274
  PIN WL275
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -480.400 -21.200 -479.400 ;
    END
  END WL275
  PIN WL276
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -482.650 -21.200 -481.650 ;
    END
  END WL276
  PIN WL277
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -484.000 -21.200 -483.000 ;
    END
  END WL277
  PIN WL278
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -486.250 -21.200 -485.250 ;
    END
  END WL278
  PIN WL279
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -487.600 -21.200 -486.600 ;
    END
  END WL279
  PIN WL280
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -489.850 -21.200 -488.850 ;
    END
  END WL280
  PIN WL281
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -491.200 -21.200 -490.200 ;
    END
  END WL281
  PIN WL282
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -493.450 -21.200 -492.450 ;
    END
  END WL282
  PIN WL283
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -494.800 -21.200 -493.800 ;
    END
  END WL283
  PIN WL284
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -497.050 -21.200 -496.050 ;
    END
  END WL284
  PIN WL285
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -498.400 -21.200 -497.400 ;
    END
  END WL285
  PIN WL286
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -500.650 -21.200 -499.650 ;
    END
  END WL286
  PIN WL287
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -502.000 -21.200 -501.000 ;
    END
  END WL287
  PIN WL288
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -504.250 -21.200 -503.250 ;
    END
  END WL288
  PIN WL289
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -505.600 -21.200 -504.600 ;
    END
  END WL289
  PIN WL290
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -507.850 -21.200 -506.850 ;
    END
  END WL290
  PIN WL291
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -509.200 -21.200 -508.200 ;
    END
  END WL291
  PIN WL292
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -511.450 -21.200 -510.450 ;
    END
  END WL292
  PIN WL293
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -512.800 -21.200 -511.800 ;
    END
  END WL293
  PIN WL294
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -515.050 -21.200 -514.050 ;
    END
  END WL294
  PIN WL295
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -516.400 -21.200 -515.400 ;
    END
  END WL295
  PIN WL296
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -518.650 -21.200 -517.650 ;
    END
  END WL296
  PIN WL297
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -520.000 -21.200 -519.000 ;
    END
  END WL297
  PIN WL298
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -522.250 -21.200 -521.250 ;
    END
  END WL298
  PIN WL299
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -523.600 -21.200 -522.600 ;
    END
  END WL299
  PIN WL300
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -525.850 -21.200 -524.850 ;
    END
  END WL300
  PIN WL301
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -527.200 -21.200 -526.200 ;
    END
  END WL301
  PIN WL302
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -529.450 -21.200 -528.450 ;
    END
  END WL302
  PIN WL303
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -530.800 -21.200 -529.800 ;
    END
  END WL303
  PIN WL304
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -533.050 -21.200 -532.050 ;
    END
  END WL304
  PIN WL305
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -534.400 -21.200 -533.400 ;
    END
  END WL305
  PIN WL306
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -536.650 -21.200 -535.650 ;
    END
  END WL306
  PIN WL307
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -538.000 -21.200 -537.000 ;
    END
  END WL307
  PIN WL308
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -540.250 -21.200 -539.250 ;
    END
  END WL308
  PIN WL309
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -541.600 -21.200 -540.600 ;
    END
  END WL309
  PIN WL310
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -543.850 -21.200 -542.850 ;
    END
  END WL310
  PIN WL311
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -545.200 -21.200 -544.200 ;
    END
  END WL311
  PIN WL312
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -547.450 -21.200 -546.450 ;
    END
  END WL312
  PIN WL313
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -548.800 -21.200 -547.800 ;
    END
  END WL313
  PIN WL314
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -551.050 -21.200 -550.050 ;
    END
  END WL314
  PIN WL315
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -552.400 -21.200 -551.400 ;
    END
  END WL315
  PIN WL316
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -554.650 -21.200 -553.650 ;
    END
  END WL316
  PIN WL317
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -556.000 -21.200 -555.000 ;
    END
  END WL317
  PIN WL318
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -558.250 -21.200 -557.250 ;
    END
  END WL318
  PIN WL319
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -559.600 -21.200 -558.600 ;
    END
  END WL319
  PIN WL320
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -561.850 -21.200 -560.850 ;
    END
  END WL320
  PIN WL321
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -563.200 -21.200 -562.200 ;
    END
  END WL321
  PIN WL322
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -565.450 -21.200 -564.450 ;
    END
  END WL322
  PIN WL323
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -566.800 -21.200 -565.800 ;
    END
  END WL323
  PIN WL324
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -569.050 -21.200 -568.050 ;
    END
  END WL324
  PIN WL325
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -570.400 -21.200 -569.400 ;
    END
  END WL325
  PIN WL326
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -572.650 -21.200 -571.650 ;
    END
  END WL326
  PIN WL327
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -574.000 -21.200 -573.000 ;
    END
  END WL327
  PIN WL328
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -576.250 -21.200 -575.250 ;
    END
  END WL328
  PIN WL329
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -577.600 -21.200 -576.600 ;
    END
  END WL329
  PIN WL330
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -579.850 -21.200 -578.850 ;
    END
  END WL330
  PIN WL331
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -581.200 -21.200 -580.200 ;
    END
  END WL331
  PIN WL332
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -583.450 -21.200 -582.450 ;
    END
  END WL332
  PIN WL333
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -584.800 -21.200 -583.800 ;
    END
  END WL333
  PIN WL334
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -587.600 -21.200 -586.600 ;
    END
  END WL334
  PIN WL335
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -588.950 -21.200 -587.950 ;
    END
  END WL335
  PIN WL336
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -591.200 -21.200 -590.200 ;
    END
  END WL336
  PIN WL337
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -592.550 -21.200 -591.550 ;
    END
  END WL337
  PIN WL338
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -594.800 -21.200 -593.800 ;
    END
  END WL338
  PIN WL339
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -596.150 -21.200 -595.150 ;
    END
  END WL339
  PIN WL340
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -598.400 -21.200 -597.400 ;
    END
  END WL340
  PIN WL341
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -599.750 -21.200 -598.750 ;
    END
  END WL341
  PIN WL342
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -602.000 -21.200 -601.000 ;
    END
  END WL342
  PIN WL343
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -603.350 -21.200 -602.350 ;
    END
  END WL343
  PIN WL344
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -605.600 -21.200 -604.600 ;
    END
  END WL344
  PIN WL345
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -606.950 -21.200 -605.950 ;
    END
  END WL345
  PIN WL346
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -609.200 -21.200 -608.200 ;
    END
  END WL346
  PIN WL347
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -610.550 -21.200 -609.550 ;
    END
  END WL347
  PIN WL348
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -612.800 -21.200 -611.800 ;
    END
  END WL348
  PIN WL349
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -614.150 -21.200 -613.150 ;
    END
  END WL349
  PIN WL350
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -616.400 -21.200 -615.400 ;
    END
  END WL350
  PIN WL351
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -617.750 -21.200 -616.750 ;
    END
  END WL351
  PIN WL352
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -620.000 -21.200 -619.000 ;
    END
  END WL352
  PIN WL353
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -621.350 -21.200 -620.350 ;
    END
  END WL353
  PIN WL354
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -623.600 -21.200 -622.600 ;
    END
  END WL354
  PIN WL355
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -624.950 -21.200 -623.950 ;
    END
  END WL355
  PIN WL356
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -627.200 -21.200 -626.200 ;
    END
  END WL356
  PIN WL357
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -628.550 -21.200 -627.550 ;
    END
  END WL357
  PIN WL358
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -630.800 -21.200 -629.800 ;
    END
  END WL358
  PIN WL359
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -632.150 -21.200 -631.150 ;
    END
  END WL359
  PIN WL360
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -634.400 -21.200 -633.400 ;
    END
  END WL360
  PIN WL361
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -635.750 -21.200 -634.750 ;
    END
  END WL361
  PIN WL362
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -638.000 -21.200 -637.000 ;
    END
  END WL362
  PIN WL363
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -639.350 -21.200 -638.350 ;
    END
  END WL363
  PIN WL364
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -641.600 -21.200 -640.600 ;
    END
  END WL364
  PIN WL365
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -642.950 -21.200 -641.950 ;
    END
  END WL365
  PIN WL366
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -645.200 -21.200 -644.200 ;
    END
  END WL366
  PIN WL367
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -646.550 -21.200 -645.550 ;
    END
  END WL367
  PIN WL368
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -648.800 -21.200 -647.800 ;
    END
  END WL368
  PIN WL369
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -650.150 -21.200 -649.150 ;
    END
  END WL369
  PIN WL370
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -652.400 -21.200 -651.400 ;
    END
  END WL370
  PIN WL371
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -653.750 -21.200 -652.750 ;
    END
  END WL371
  PIN WL372
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -656.000 -21.200 -655.000 ;
    END
  END WL372
  PIN WL373
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -657.350 -21.200 -656.350 ;
    END
  END WL373
  PIN WL374
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -659.600 -21.200 -658.600 ;
    END
  END WL374
  PIN WL375
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -660.950 -21.200 -659.950 ;
    END
  END WL375
  PIN WL376
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -663.200 -21.200 -662.200 ;
    END
  END WL376
  PIN WL377
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -664.550 -21.200 -663.550 ;
    END
  END WL377
  PIN WL378
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -666.800 -21.200 -665.800 ;
    END
  END WL378
  PIN WL379
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -668.150 -21.200 -667.150 ;
    END
  END WL379
  PIN WL380
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -670.400 -21.200 -669.400 ;
    END
  END WL380
  PIN WL381
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -671.750 -21.200 -670.750 ;
    END
  END WL381
  PIN WL382
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -674.000 -21.200 -673.000 ;
    END
  END WL382
  PIN WL383
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -675.350 -21.200 -674.350 ;
    END
  END WL383
  PIN WL384
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -677.600 -21.200 -676.600 ;
    END
  END WL384
  PIN WL385
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -678.950 -21.200 -677.950 ;
    END
  END WL385
  PIN WL386
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -681.200 -21.200 -680.200 ;
    END
  END WL386
  PIN WL387
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -682.550 -21.200 -681.550 ;
    END
  END WL387
  PIN WL388
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -684.800 -21.200 -683.800 ;
    END
  END WL388
  PIN WL389
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -686.150 -21.200 -685.150 ;
    END
  END WL389
  PIN WL390
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -688.400 -21.200 -687.400 ;
    END
  END WL390
  PIN WL391
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -689.750 -21.200 -688.750 ;
    END
  END WL391
  PIN WL392
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -692.000 -21.200 -691.000 ;
    END
  END WL392
  PIN WL393
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -693.350 -21.200 -692.350 ;
    END
  END WL393
  PIN WL394
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -695.600 -21.200 -694.600 ;
    END
  END WL394
  PIN WL395
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -696.950 -21.200 -695.950 ;
    END
  END WL395
  PIN WL396
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -699.200 -21.200 -698.200 ;
    END
  END WL396
  PIN WL397
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -700.550 -21.200 -699.550 ;
    END
  END WL397
  PIN WL398
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -702.800 -21.200 -701.800 ;
    END
  END WL398
  PIN WL399
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -704.150 -21.200 -703.150 ;
    END
  END WL399
  PIN WL400
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -706.400 -21.200 -705.400 ;
    END
  END WL400
  PIN WL401
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -707.750 -21.200 -706.750 ;
    END
  END WL401
  PIN WL402
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -710.000 -21.200 -709.000 ;
    END
  END WL402
  PIN WL403
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -711.350 -21.200 -710.350 ;
    END
  END WL403
  PIN WL404
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -713.600 -21.200 -712.600 ;
    END
  END WL404
  PIN WL405
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -714.950 -21.200 -713.950 ;
    END
  END WL405
  PIN WL406
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -717.200 -21.200 -716.200 ;
    END
  END WL406
  PIN WL407
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -718.550 -21.200 -717.550 ;
    END
  END WL407
  PIN WL408
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -720.800 -21.200 -719.800 ;
    END
  END WL408
  PIN WL409
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -722.150 -21.200 -721.150 ;
    END
  END WL409
  PIN WL410
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -724.400 -21.200 -723.400 ;
    END
  END WL410
  PIN WL411
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -725.750 -21.200 -724.750 ;
    END
  END WL411
  PIN WL412
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -728.000 -21.200 -727.000 ;
    END
  END WL412
  PIN WL413
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -729.350 -21.200 -728.350 ;
    END
  END WL413
  PIN WL414
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -731.600 -21.200 -730.600 ;
    END
  END WL414
  PIN WL415
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -732.950 -21.200 -731.950 ;
    END
  END WL415
  PIN WL416
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -735.200 -21.200 -734.200 ;
    END
  END WL416
  PIN WL417
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -736.550 -21.200 -735.550 ;
    END
  END WL417
  PIN WL418
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -738.800 -21.200 -737.800 ;
    END
  END WL418
  PIN WL419
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -740.150 -21.200 -739.150 ;
    END
  END WL419
  PIN WL420
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -742.400 -21.200 -741.400 ;
    END
  END WL420
  PIN WL421
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -743.750 -21.200 -742.750 ;
    END
  END WL421
  PIN WL422
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -746.000 -21.200 -745.000 ;
    END
  END WL422
  PIN WL423
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -747.350 -21.200 -746.350 ;
    END
  END WL423
  PIN WL424
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -749.600 -21.200 -748.600 ;
    END
  END WL424
  PIN WL425
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -750.950 -21.200 -749.950 ;
    END
  END WL425
  PIN WL426
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -753.200 -21.200 -752.200 ;
    END
  END WL426
  PIN WL427
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -754.550 -21.200 -753.550 ;
    END
  END WL427
  PIN WL428
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -756.800 -21.200 -755.800 ;
    END
  END WL428
  PIN WL429
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -758.150 -21.200 -757.150 ;
    END
  END WL429
  PIN WL430
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -760.400 -21.200 -759.400 ;
    END
  END WL430
  PIN WL431
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -761.750 -21.200 -760.750 ;
    END
  END WL431
  PIN WL432
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -764.000 -21.200 -763.000 ;
    END
  END WL432
  PIN WL433
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -765.350 -21.200 -764.350 ;
    END
  END WL433
  PIN WL434
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -767.600 -21.200 -766.600 ;
    END
  END WL434
  PIN WL435
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -768.950 -21.200 -767.950 ;
    END
  END WL435
  PIN WL436
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -771.200 -21.200 -770.200 ;
    END
  END WL436
  PIN WL437
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -772.550 -21.200 -771.550 ;
    END
  END WL437
  PIN WL438
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -774.800 -21.200 -773.800 ;
    END
  END WL438
  PIN WL439
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -776.150 -21.200 -775.150 ;
    END
  END WL439
  PIN WL440
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -778.400 -21.200 -777.400 ;
    END
  END WL440
  PIN WL441
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -779.750 -21.200 -778.750 ;
    END
  END WL441
  PIN WL442
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -782.000 -21.200 -781.000 ;
    END
  END WL442
  PIN WL443
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -783.350 -21.200 -782.350 ;
    END
  END WL443
  PIN WL444
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -786.150 -21.200 -785.150 ;
    END
  END WL444
  PIN WL445
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -787.500 -21.200 -786.500 ;
    END
  END WL445
  PIN WL446
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -789.750 -21.200 -788.750 ;
    END
  END WL446
  PIN WL447
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -791.100 -21.200 -790.100 ;
    END
  END WL447
  PIN WL448
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -793.350 -21.200 -792.350 ;
    END
  END WL448
  PIN WL449
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -794.700 -21.200 -793.700 ;
    END
  END WL449
  PIN WL450
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -796.950 -21.200 -795.950 ;
    END
  END WL450
  PIN WL451
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -798.300 -21.200 -797.300 ;
    END
  END WL451
  PIN WL452
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -800.550 -21.200 -799.550 ;
    END
  END WL452
  PIN WL453
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -801.900 -21.200 -800.900 ;
    END
  END WL453
  PIN WL454
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -804.150 -21.200 -803.150 ;
    END
  END WL454
  PIN WL455
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -805.500 -21.200 -804.500 ;
    END
  END WL455
  PIN WL456
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -807.750 -21.200 -806.750 ;
    END
  END WL456
  PIN WL457
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -809.100 -21.200 -808.100 ;
    END
  END WL457
  PIN WL458
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -811.350 -21.200 -810.350 ;
    END
  END WL458
  PIN WL459
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -812.700 -21.200 -811.700 ;
    END
  END WL459
  PIN WL460
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -814.950 -21.200 -813.950 ;
    END
  END WL460
  PIN WL461
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -816.300 -21.200 -815.300 ;
    END
  END WL461
  PIN WL462
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -818.550 -21.200 -817.550 ;
    END
  END WL462
  PIN WL463
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -819.900 -21.200 -818.900 ;
    END
  END WL463
  PIN WL464
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -822.150 -21.200 -821.150 ;
    END
  END WL464
  PIN WL465
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -823.500 -21.200 -822.500 ;
    END
  END WL465
  PIN WL466
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -825.750 -21.200 -824.750 ;
    END
  END WL466
  PIN WL467
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -827.100 -21.200 -826.100 ;
    END
  END WL467
  PIN WL468
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -829.350 -21.200 -828.350 ;
    END
  END WL468
  PIN WL469
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -830.700 -21.200 -829.700 ;
    END
  END WL469
  PIN WL470
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -832.950 -21.200 -831.950 ;
    END
  END WL470
  PIN WL471
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -834.300 -21.200 -833.300 ;
    END
  END WL471
  PIN WL472
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -836.550 -21.200 -835.550 ;
    END
  END WL472
  PIN WL473
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -837.900 -21.200 -836.900 ;
    END
  END WL473
  PIN WL474
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -840.150 -21.200 -839.150 ;
    END
  END WL474
  PIN WL475
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -841.500 -21.200 -840.500 ;
    END
  END WL475
  PIN WL476
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -843.750 -21.200 -842.750 ;
    END
  END WL476
  PIN WL477
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -845.100 -21.200 -844.100 ;
    END
  END WL477
  PIN WL478
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -847.350 -21.200 -846.350 ;
    END
  END WL478
  PIN WL479
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -848.700 -21.200 -847.700 ;
    END
  END WL479
  PIN WL480
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -850.950 -21.200 -849.950 ;
    END
  END WL480
  PIN WL481
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -852.300 -21.200 -851.300 ;
    END
  END WL481
  PIN WL482
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -854.550 -21.200 -853.550 ;
    END
  END WL482
  PIN WL483
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -855.900 -21.200 -854.900 ;
    END
  END WL483
  PIN WL484
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -858.150 -21.200 -857.150 ;
    END
  END WL484
  PIN WL485
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -859.500 -21.200 -858.500 ;
    END
  END WL485
  PIN WL486
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -861.750 -21.200 -860.750 ;
    END
  END WL486
  PIN WL487
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -863.100 -21.200 -862.100 ;
    END
  END WL487
  PIN WL488
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -865.350 -21.200 -864.350 ;
    END
  END WL488
  PIN WL489
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -866.700 -21.200 -865.700 ;
    END
  END WL489
  PIN WL490
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -868.950 -21.200 -867.950 ;
    END
  END WL490
  PIN WL491
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -870.300 -21.200 -869.300 ;
    END
  END WL491
  PIN WL492
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -872.550 -21.200 -871.550 ;
    END
  END WL492
  PIN WL493
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -873.900 -21.200 -872.900 ;
    END
  END WL493
  PIN WL494
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -876.150 -21.200 -875.150 ;
    END
  END WL494
  PIN WL495
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -877.500 -21.200 -876.500 ;
    END
  END WL495
  PIN WL496
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -879.750 -21.200 -878.750 ;
    END
  END WL496
  PIN WL497
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -881.100 -21.200 -880.100 ;
    END
  END WL497
  PIN WL498
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -883.350 -21.200 -882.350 ;
    END
  END WL498
  PIN WL499
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -884.700 -21.200 -883.700 ;
    END
  END WL499
  PIN WL500
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -886.950 -21.200 -885.950 ;
    END
  END WL500
  PIN WL501
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -888.300 -21.200 -887.300 ;
    END
  END WL501
  PIN WL502
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -890.550 -21.200 -889.550 ;
    END
  END WL502
  PIN WL503
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -891.900 -21.200 -890.900 ;
    END
  END WL503
  PIN WL504
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -894.150 -21.200 -893.150 ;
    END
  END WL504
  PIN WL505
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -895.500 -21.200 -894.500 ;
    END
  END WL505
  PIN WL506
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -897.750 -21.200 -896.750 ;
    END
  END WL506
  PIN WL507
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -899.100 -21.200 -898.100 ;
    END
  END WL507
  PIN WL508
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -901.350 -21.200 -900.350 ;
    END
  END WL508
  PIN WL509
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -902.700 -21.200 -901.700 ;
    END
  END WL509
  PIN WL510
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -904.950 -21.200 -903.950 ;
    END
  END WL510
  PIN WL511
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -906.300 -21.200 -905.300 ;
    END
  END WL511
  PIN WL512
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -908.550 -21.200 -907.550 ;
    END
  END WL512
  PIN WL513
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -909.900 -21.200 -908.900 ;
    END
  END WL513
  PIN WL514
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -912.150 -21.200 -911.150 ;
    END
  END WL514
  PIN WL515
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -913.500 -21.200 -912.500 ;
    END
  END WL515
  PIN WL516
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -915.750 -21.200 -914.750 ;
    END
  END WL516
  PIN WL517
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -917.100 -21.200 -916.100 ;
    END
  END WL517
  PIN WL518
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -919.350 -21.200 -918.350 ;
    END
  END WL518
  PIN WL519
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -920.700 -21.200 -919.700 ;
    END
  END WL519
  PIN WL520
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -922.950 -21.200 -921.950 ;
    END
  END WL520
  PIN WL521
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -924.300 -21.200 -923.300 ;
    END
  END WL521
  PIN WL522
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -926.550 -21.200 -925.550 ;
    END
  END WL522
  PIN WL523
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -927.900 -21.200 -926.900 ;
    END
  END WL523
  PIN WL524
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -930.150 -21.200 -929.150 ;
    END
  END WL524
  PIN WL525
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -931.500 -21.200 -930.500 ;
    END
  END WL525
  PIN WL526
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -933.750 -21.200 -932.750 ;
    END
  END WL526
  PIN WL527
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -935.100 -21.200 -934.100 ;
    END
  END WL527
  PIN WL528
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -937.350 -21.200 -936.350 ;
    END
  END WL528
  PIN WL529
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -938.700 -21.200 -937.700 ;
    END
  END WL529
  PIN WL530
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -940.950 -21.200 -939.950 ;
    END
  END WL530
  PIN WL531
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -942.300 -21.200 -941.300 ;
    END
  END WL531
  PIN WL532
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -944.550 -21.200 -943.550 ;
    END
  END WL532
  PIN WL533
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -945.900 -21.200 -944.900 ;
    END
  END WL533
  PIN WL534
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -948.150 -21.200 -947.150 ;
    END
  END WL534
  PIN WL535
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -949.500 -21.200 -948.500 ;
    END
  END WL535
  PIN WL536
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -951.750 -21.200 -950.750 ;
    END
  END WL536
  PIN WL537
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -953.100 -21.200 -952.100 ;
    END
  END WL537
  PIN WL538
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -955.350 -21.200 -954.350 ;
    END
  END WL538
  PIN WL539
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -956.700 -21.200 -955.700 ;
    END
  END WL539
  PIN WL540
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -958.950 -21.200 -957.950 ;
    END
  END WL540
  PIN WL541
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -960.300 -21.200 -959.300 ;
    END
  END WL541
  PIN WL542
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -962.550 -21.200 -961.550 ;
    END
  END WL542
  PIN WL543
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -963.900 -21.200 -962.900 ;
    END
  END WL543
  PIN WL544
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -966.150 -21.200 -965.150 ;
    END
  END WL544
  PIN WL545
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -967.500 -21.200 -966.500 ;
    END
  END WL545
  PIN WL546
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -969.750 -21.200 -968.750 ;
    END
  END WL546
  PIN WL547
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -971.100 -21.200 -970.100 ;
    END
  END WL547
  PIN WL548
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -973.350 -21.200 -972.350 ;
    END
  END WL548
  PIN WL549
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -974.700 -21.200 -973.700 ;
    END
  END WL549
  PIN WL550
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -976.950 -21.200 -975.950 ;
    END
  END WL550
  PIN WL551
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -978.300 -21.200 -977.300 ;
    END
  END WL551
  PIN WL552
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -980.550 -21.200 -979.550 ;
    END
  END WL552
  PIN WL553
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -981.900 -21.200 -980.900 ;
    END
  END WL553
  PIN WL554
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -984.700 -21.200 -983.700 ;
    END
  END WL554
  PIN WL555
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -986.050 -21.200 -985.050 ;
    END
  END WL555
  PIN WL556
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -988.300 -21.200 -987.300 ;
    END
  END WL556
  PIN WL557
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -989.650 -21.200 -988.650 ;
    END
  END WL557
  PIN WL558
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -991.900 -21.200 -990.900 ;
    END
  END WL558
  PIN WL559
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -993.250 -21.200 -992.250 ;
    END
  END WL559
  PIN WL560
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -995.500 -21.200 -994.500 ;
    END
  END WL560
  PIN WL561
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -996.850 -21.200 -995.850 ;
    END
  END WL561
  PIN WL562
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -999.100 -21.200 -998.100 ;
    END
  END WL562
  PIN WL563
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1000.450 -21.200 -999.450 ;
    END
  END WL563
  PIN WL564
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1002.700 -21.200 -1001.700 ;
    END
  END WL564
  PIN WL565
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1004.050 -21.200 -1003.050 ;
    END
  END WL565
  PIN WL566
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1006.300 -21.200 -1005.300 ;
    END
  END WL566
  PIN WL567
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1007.650 -21.200 -1006.650 ;
    END
  END WL567
  PIN WL568
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1009.900 -21.200 -1008.900 ;
    END
  END WL568
  PIN WL569
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1011.250 -21.200 -1010.250 ;
    END
  END WL569
  PIN WL570
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1013.500 -21.200 -1012.500 ;
    END
  END WL570
  PIN WL571
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1014.850 -21.200 -1013.850 ;
    END
  END WL571
  PIN WL572
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1017.100 -21.200 -1016.100 ;
    END
  END WL572
  PIN WL573
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1018.450 -21.200 -1017.450 ;
    END
  END WL573
  PIN WL574
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1020.700 -21.200 -1019.700 ;
    END
  END WL574
  PIN WL575
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1022.050 -21.200 -1021.050 ;
    END
  END WL575
  PIN WL576
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1024.300 -21.200 -1023.300 ;
    END
  END WL576
  PIN WL577
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1025.650 -21.200 -1024.650 ;
    END
  END WL577
  PIN WL578
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1027.900 -21.200 -1026.900 ;
    END
  END WL578
  PIN WL579
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1029.250 -21.200 -1028.250 ;
    END
  END WL579
  PIN WL580
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1031.500 -21.200 -1030.500 ;
    END
  END WL580
  PIN WL581
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1032.850 -21.200 -1031.850 ;
    END
  END WL581
  PIN WL582
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1035.100 -21.200 -1034.100 ;
    END
  END WL582
  PIN WL583
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1036.450 -21.200 -1035.450 ;
    END
  END WL583
  PIN WL584
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1038.700 -21.200 -1037.700 ;
    END
  END WL584
  PIN WL585
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1040.050 -21.200 -1039.050 ;
    END
  END WL585
  PIN WL586
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1042.300 -21.200 -1041.300 ;
    END
  END WL586
  PIN WL587
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1043.650 -21.200 -1042.650 ;
    END
  END WL587
  PIN WL588
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1045.900 -21.200 -1044.900 ;
    END
  END WL588
  PIN WL589
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1047.250 -21.200 -1046.250 ;
    END
  END WL589
  PIN WL590
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1049.500 -21.200 -1048.500 ;
    END
  END WL590
  PIN WL591
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1050.850 -21.200 -1049.850 ;
    END
  END WL591
  PIN WL592
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1053.100 -21.200 -1052.100 ;
    END
  END WL592
  PIN WL593
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1054.450 -21.200 -1053.450 ;
    END
  END WL593
  PIN WL594
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1056.700 -21.200 -1055.700 ;
    END
  END WL594
  PIN WL595
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1058.050 -21.200 -1057.050 ;
    END
  END WL595
  PIN WL596
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1060.300 -21.200 -1059.300 ;
    END
  END WL596
  PIN WL597
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1061.650 -21.200 -1060.650 ;
    END
  END WL597
  PIN WL598
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1063.900 -21.200 -1062.900 ;
    END
  END WL598
  PIN WL599
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1065.250 -21.200 -1064.250 ;
    END
  END WL599
  PIN WL600
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1067.500 -21.200 -1066.500 ;
    END
  END WL600
  PIN WL601
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1068.850 -21.200 -1067.850 ;
    END
  END WL601
  PIN WL602
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1071.100 -21.200 -1070.100 ;
    END
  END WL602
  PIN WL603
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1072.450 -21.200 -1071.450 ;
    END
  END WL603
  PIN WL604
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1074.700 -21.200 -1073.700 ;
    END
  END WL604
  PIN WL605
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1076.050 -21.200 -1075.050 ;
    END
  END WL605
  PIN WL606
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1078.300 -21.200 -1077.300 ;
    END
  END WL606
  PIN WL607
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1079.650 -21.200 -1078.650 ;
    END
  END WL607
  PIN WL608
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1081.900 -21.200 -1080.900 ;
    END
  END WL608
  PIN WL609
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1083.250 -21.200 -1082.250 ;
    END
  END WL609
  PIN WL610
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1085.500 -21.200 -1084.500 ;
    END
  END WL610
  PIN WL611
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1086.850 -21.200 -1085.850 ;
    END
  END WL611
  PIN WL612
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1089.100 -21.200 -1088.100 ;
    END
  END WL612
  PIN WL613
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1090.450 -21.200 -1089.450 ;
    END
  END WL613
  PIN WL614
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1092.700 -21.200 -1091.700 ;
    END
  END WL614
  PIN WL615
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1094.050 -21.200 -1093.050 ;
    END
  END WL615
  PIN WL616
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1096.300 -21.200 -1095.300 ;
    END
  END WL616
  PIN WL617
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1097.650 -21.200 -1096.650 ;
    END
  END WL617
  PIN WL618
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1099.900 -21.200 -1098.900 ;
    END
  END WL618
  PIN WL619
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1101.250 -21.200 -1100.250 ;
    END
  END WL619
  PIN WL620
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1103.500 -21.200 -1102.500 ;
    END
  END WL620
  PIN WL621
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1104.850 -21.200 -1103.850 ;
    END
  END WL621
  PIN WL622
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1107.100 -21.200 -1106.100 ;
    END
  END WL622
  PIN WL623
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1108.450 -21.200 -1107.450 ;
    END
  END WL623
  PIN WL624
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1110.700 -21.200 -1109.700 ;
    END
  END WL624
  PIN WL625
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1112.050 -21.200 -1111.050 ;
    END
  END WL625
  PIN WL626
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1114.300 -21.200 -1113.300 ;
    END
  END WL626
  PIN WL627
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1115.650 -21.200 -1114.650 ;
    END
  END WL627
  PIN WL628
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1117.900 -21.200 -1116.900 ;
    END
  END WL628
  PIN WL629
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1119.250 -21.200 -1118.250 ;
    END
  END WL629
  PIN WL630
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1121.500 -21.200 -1120.500 ;
    END
  END WL630
  PIN WL631
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1122.850 -21.200 -1121.850 ;
    END
  END WL631
  PIN WL632
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1125.100 -21.200 -1124.100 ;
    END
  END WL632
  PIN WL633
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1126.450 -21.200 -1125.450 ;
    END
  END WL633
  PIN WL634
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1128.700 -21.200 -1127.700 ;
    END
  END WL634
  PIN WL635
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1130.050 -21.200 -1129.050 ;
    END
  END WL635
  PIN WL636
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1132.300 -21.200 -1131.300 ;
    END
  END WL636
  PIN WL637
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1133.650 -21.200 -1132.650 ;
    END
  END WL637
  PIN WL638
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1135.900 -21.200 -1134.900 ;
    END
  END WL638
  PIN WL639
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1137.250 -21.200 -1136.250 ;
    END
  END WL639
  PIN WL640
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1139.500 -21.200 -1138.500 ;
    END
  END WL640
  PIN WL641
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1140.850 -21.200 -1139.850 ;
    END
  END WL641
  PIN WL642
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1143.100 -21.200 -1142.100 ;
    END
  END WL642
  PIN WL643
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1144.450 -21.200 -1143.450 ;
    END
  END WL643
  PIN WL644
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1146.700 -21.200 -1145.700 ;
    END
  END WL644
  PIN WL645
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1148.050 -21.200 -1147.050 ;
    END
  END WL645
  PIN WL646
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1150.300 -21.200 -1149.300 ;
    END
  END WL646
  PIN WL647
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1151.650 -21.200 -1150.650 ;
    END
  END WL647
  PIN WL648
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1153.900 -21.200 -1152.900 ;
    END
  END WL648
  PIN WL649
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1155.250 -21.200 -1154.250 ;
    END
  END WL649
  PIN WL650
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1157.500 -21.200 -1156.500 ;
    END
  END WL650
  PIN WL651
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1158.850 -21.200 -1157.850 ;
    END
  END WL651
  PIN WL652
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1161.100 -21.200 -1160.100 ;
    END
  END WL652
  PIN WL653
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1162.450 -21.200 -1161.450 ;
    END
  END WL653
  PIN WL654
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1164.700 -21.200 -1163.700 ;
    END
  END WL654
  PIN WL655
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1166.050 -21.200 -1165.050 ;
    END
  END WL655
  PIN WL656
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1168.300 -21.200 -1167.300 ;
    END
  END WL656
  PIN WL657
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1169.650 -21.200 -1168.650 ;
    END
  END WL657
  PIN WL658
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1171.900 -21.200 -1170.900 ;
    END
  END WL658
  PIN WL659
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1173.250 -21.200 -1172.250 ;
    END
  END WL659
  PIN WL660
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1175.500 -21.200 -1174.500 ;
    END
  END WL660
  PIN WL661
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1176.850 -21.200 -1175.850 ;
    END
  END WL661
  PIN WL662
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1179.100 -21.200 -1178.100 ;
    END
  END WL662
  PIN WL663
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1180.450 -21.200 -1179.450 ;
    END
  END WL663
  PIN WL664
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1183.250 -21.200 -1182.250 ;
    END
  END WL664
  PIN WL665
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1184.600 -21.200 -1183.600 ;
    END
  END WL665
  PIN WL666
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1186.850 -21.200 -1185.850 ;
    END
  END WL666
  PIN WL667
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1188.200 -21.200 -1187.200 ;
    END
  END WL667
  PIN WL668
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1190.450 -21.200 -1189.450 ;
    END
  END WL668
  PIN WL669
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1191.800 -21.200 -1190.800 ;
    END
  END WL669
  PIN WL670
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1194.050 -21.200 -1193.050 ;
    END
  END WL670
  PIN WL671
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1195.400 -21.200 -1194.400 ;
    END
  END WL671
  PIN WL672
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1197.650 -21.200 -1196.650 ;
    END
  END WL672
  PIN WL673
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1199.000 -21.200 -1198.000 ;
    END
  END WL673
  PIN WL674
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1201.250 -21.200 -1200.250 ;
    END
  END WL674
  PIN WL675
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1202.600 -21.200 -1201.600 ;
    END
  END WL675
  PIN WL676
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1204.850 -21.200 -1203.850 ;
    END
  END WL676
  PIN WL677
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1206.200 -21.200 -1205.200 ;
    END
  END WL677
  PIN WL678
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1208.450 -21.200 -1207.450 ;
    END
  END WL678
  PIN WL679
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1209.800 -21.200 -1208.800 ;
    END
  END WL679
  PIN WL680
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1212.050 -21.200 -1211.050 ;
    END
  END WL680
  PIN WL681
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1213.400 -21.200 -1212.400 ;
    END
  END WL681
  PIN WL682
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1215.650 -21.200 -1214.650 ;
    END
  END WL682
  PIN WL683
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1217.000 -21.200 -1216.000 ;
    END
  END WL683
  PIN WL684
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1219.250 -21.200 -1218.250 ;
    END
  END WL684
  PIN WL685
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1220.600 -21.200 -1219.600 ;
    END
  END WL685
  PIN WL686
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1222.850 -21.200 -1221.850 ;
    END
  END WL686
  PIN WL687
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1224.200 -21.200 -1223.200 ;
    END
  END WL687
  PIN WL688
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1226.450 -21.200 -1225.450 ;
    END
  END WL688
  PIN WL689
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1227.800 -21.200 -1226.800 ;
    END
  END WL689
  PIN WL690
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1230.050 -21.200 -1229.050 ;
    END
  END WL690
  PIN WL691
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1231.400 -21.200 -1230.400 ;
    END
  END WL691
  PIN WL692
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1233.650 -21.200 -1232.650 ;
    END
  END WL692
  PIN WL693
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1235.000 -21.200 -1234.000 ;
    END
  END WL693
  PIN WL694
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1237.250 -21.200 -1236.250 ;
    END
  END WL694
  PIN WL695
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1238.600 -21.200 -1237.600 ;
    END
  END WL695
  PIN WL696
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1240.850 -21.200 -1239.850 ;
    END
  END WL696
  PIN WL697
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1242.200 -21.200 -1241.200 ;
    END
  END WL697
  PIN WL698
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1244.450 -21.200 -1243.450 ;
    END
  END WL698
  PIN WL699
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1245.800 -21.200 -1244.800 ;
    END
  END WL699
  PIN WL700
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1248.050 -21.200 -1247.050 ;
    END
  END WL700
  PIN WL701
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1249.400 -21.200 -1248.400 ;
    END
  END WL701
  PIN WL702
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1251.650 -21.200 -1250.650 ;
    END
  END WL702
  PIN WL703
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1253.000 -21.200 -1252.000 ;
    END
  END WL703
  PIN WL704
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1255.250 -21.200 -1254.250 ;
    END
  END WL704
  PIN WL705
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1256.600 -21.200 -1255.600 ;
    END
  END WL705
  PIN WL706
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1258.850 -21.200 -1257.850 ;
    END
  END WL706
  PIN WL707
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1260.200 -21.200 -1259.200 ;
    END
  END WL707
  PIN WL708
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1262.450 -21.200 -1261.450 ;
    END
  END WL708
  PIN WL709
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1263.800 -21.200 -1262.800 ;
    END
  END WL709
  PIN WL710
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1266.050 -21.200 -1265.050 ;
    END
  END WL710
  PIN WL711
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1267.400 -21.200 -1266.400 ;
    END
  END WL711
  PIN WL712
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1269.650 -21.200 -1268.650 ;
    END
  END WL712
  PIN WL713
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1271.000 -21.200 -1270.000 ;
    END
  END WL713
  PIN WL714
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1273.250 -21.200 -1272.250 ;
    END
  END WL714
  PIN WL715
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1274.600 -21.200 -1273.600 ;
    END
  END WL715
  PIN WL716
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1276.850 -21.200 -1275.850 ;
    END
  END WL716
  PIN WL717
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1278.200 -21.200 -1277.200 ;
    END
  END WL717
  PIN WL718
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1280.450 -21.200 -1279.450 ;
    END
  END WL718
  PIN WL719
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1281.800 -21.200 -1280.800 ;
    END
  END WL719
  PIN WL720
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1284.050 -21.200 -1283.050 ;
    END
  END WL720
  PIN WL721
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1285.400 -21.200 -1284.400 ;
    END
  END WL721
  PIN WL722
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1287.650 -21.200 -1286.650 ;
    END
  END WL722
  PIN WL723
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1289.000 -21.200 -1288.000 ;
    END
  END WL723
  PIN WL724
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1291.250 -21.200 -1290.250 ;
    END
  END WL724
  PIN WL725
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1292.600 -21.200 -1291.600 ;
    END
  END WL725
  PIN WL726
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1294.850 -21.200 -1293.850 ;
    END
  END WL726
  PIN WL727
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1296.200 -21.200 -1295.200 ;
    END
  END WL727
  PIN WL728
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1298.450 -21.200 -1297.450 ;
    END
  END WL728
  PIN WL729
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1299.800 -21.200 -1298.800 ;
    END
  END WL729
  PIN WL730
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1302.050 -21.200 -1301.050 ;
    END
  END WL730
  PIN WL731
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1303.400 -21.200 -1302.400 ;
    END
  END WL731
  PIN WL732
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1305.650 -21.200 -1304.650 ;
    END
  END WL732
  PIN WL733
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1307.000 -21.200 -1306.000 ;
    END
  END WL733
  PIN WL734
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1309.250 -21.200 -1308.250 ;
    END
  END WL734
  PIN WL735
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1310.600 -21.200 -1309.600 ;
    END
  END WL735
  PIN WL736
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1312.850 -21.200 -1311.850 ;
    END
  END WL736
  PIN WL737
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1314.200 -21.200 -1313.200 ;
    END
  END WL737
  PIN WL738
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1316.450 -21.200 -1315.450 ;
    END
  END WL738
  PIN WL739
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1317.800 -21.200 -1316.800 ;
    END
  END WL739
  PIN WL740
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1320.050 -21.200 -1319.050 ;
    END
  END WL740
  PIN WL741
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1321.400 -21.200 -1320.400 ;
    END
  END WL741
  PIN WL742
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1323.650 -21.200 -1322.650 ;
    END
  END WL742
  PIN WL743
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1325.000 -21.200 -1324.000 ;
    END
  END WL743
  PIN WL744
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1327.250 -21.200 -1326.250 ;
    END
  END WL744
  PIN WL745
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1328.600 -21.200 -1327.600 ;
    END
  END WL745
  PIN WL746
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1330.850 -21.200 -1329.850 ;
    END
  END WL746
  PIN WL747
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1332.200 -21.200 -1331.200 ;
    END
  END WL747
  PIN WL748
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1334.450 -21.200 -1333.450 ;
    END
  END WL748
  PIN WL749
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1335.800 -21.200 -1334.800 ;
    END
  END WL749
  PIN WL750
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1338.050 -21.200 -1337.050 ;
    END
  END WL750
  PIN WL751
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1339.400 -21.200 -1338.400 ;
    END
  END WL751
  PIN WL752
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1341.650 -21.200 -1340.650 ;
    END
  END WL752
  PIN WL753
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1343.000 -21.200 -1342.000 ;
    END
  END WL753
  PIN WL754
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1345.250 -21.200 -1344.250 ;
    END
  END WL754
  PIN WL755
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1346.600 -21.200 -1345.600 ;
    END
  END WL755
  PIN WL756
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1348.850 -21.200 -1347.850 ;
    END
  END WL756
  PIN WL757
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1350.200 -21.200 -1349.200 ;
    END
  END WL757
  PIN WL758
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1352.450 -21.200 -1351.450 ;
    END
  END WL758
  PIN WL759
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1353.800 -21.200 -1352.800 ;
    END
  END WL759
  PIN WL760
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1356.050 -21.200 -1355.050 ;
    END
  END WL760
  PIN WL761
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1357.400 -21.200 -1356.400 ;
    END
  END WL761
  PIN WL762
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1359.650 -21.200 -1358.650 ;
    END
  END WL762
  PIN WL763
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1361.000 -21.200 -1360.000 ;
    END
  END WL763
  PIN WL764
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1363.250 -21.200 -1362.250 ;
    END
  END WL764
  PIN WL765
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1364.600 -21.200 -1363.600 ;
    END
  END WL765
  PIN WL766
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1366.850 -21.200 -1365.850 ;
    END
  END WL766
  PIN WL767
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1368.200 -21.200 -1367.200 ;
    END
  END WL767
  PIN WL768
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1370.450 -21.200 -1369.450 ;
    END
  END WL768
  PIN WL769
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1371.800 -21.200 -1370.800 ;
    END
  END WL769
  PIN WL770
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1374.050 -21.200 -1373.050 ;
    END
  END WL770
  PIN WL771
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1375.400 -21.200 -1374.400 ;
    END
  END WL771
  PIN WL772
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1377.650 -21.200 -1376.650 ;
    END
  END WL772
  PIN WL773
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1379.000 -21.200 -1378.000 ;
    END
  END WL773
  PIN WL774
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1381.800 -21.200 -1380.800 ;
    END
  END WL774
  PIN WL775
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1383.150 -21.200 -1382.150 ;
    END
  END WL775
  PIN WL776
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1385.400 -21.200 -1384.400 ;
    END
  END WL776
  PIN WL777
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1386.750 -21.200 -1385.750 ;
    END
  END WL777
  PIN WL778
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1389.000 -21.200 -1388.000 ;
    END
  END WL778
  PIN WL779
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1390.350 -21.200 -1389.350 ;
    END
  END WL779
  PIN WL780
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1392.600 -21.200 -1391.600 ;
    END
  END WL780
  PIN WL781
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1393.950 -21.200 -1392.950 ;
    END
  END WL781
  PIN WL782
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1396.200 -21.200 -1395.200 ;
    END
  END WL782
  PIN WL783
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1397.550 -21.200 -1396.550 ;
    END
  END WL783
  PIN WL784
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1399.800 -21.200 -1398.800 ;
    END
  END WL784
  PIN WL785
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1401.150 -21.200 -1400.150 ;
    END
  END WL785
  PIN WL786
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1403.400 -21.200 -1402.400 ;
    END
  END WL786
  PIN WL787
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1404.750 -21.200 -1403.750 ;
    END
  END WL787
  PIN WL788
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1407.000 -21.200 -1406.000 ;
    END
  END WL788
  PIN WL789
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1408.350 -21.200 -1407.350 ;
    END
  END WL789
  PIN WL790
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1410.600 -21.200 -1409.600 ;
    END
  END WL790
  PIN WL791
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1411.950 -21.200 -1410.950 ;
    END
  END WL791
  PIN WL792
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1414.200 -21.200 -1413.200 ;
    END
  END WL792
  PIN WL793
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1415.550 -21.200 -1414.550 ;
    END
  END WL793
  PIN WL794
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1417.800 -21.200 -1416.800 ;
    END
  END WL794
  PIN WL795
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1419.150 -21.200 -1418.150 ;
    END
  END WL795
  PIN WL796
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1421.400 -21.200 -1420.400 ;
    END
  END WL796
  PIN WL797
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1422.750 -21.200 -1421.750 ;
    END
  END WL797
  PIN WL798
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1425.000 -21.200 -1424.000 ;
    END
  END WL798
  PIN WL799
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1426.350 -21.200 -1425.350 ;
    END
  END WL799
  PIN WL800
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1428.600 -21.200 -1427.600 ;
    END
  END WL800
  PIN WL801
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1429.950 -21.200 -1428.950 ;
    END
  END WL801
  PIN WL802
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1432.200 -21.200 -1431.200 ;
    END
  END WL802
  PIN WL803
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1433.550 -21.200 -1432.550 ;
    END
  END WL803
  PIN WL804
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1435.800 -21.200 -1434.800 ;
    END
  END WL804
  PIN WL805
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1437.150 -21.200 -1436.150 ;
    END
  END WL805
  PIN WL806
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1439.400 -21.200 -1438.400 ;
    END
  END WL806
  PIN WL807
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1440.750 -21.200 -1439.750 ;
    END
  END WL807
  PIN WL808
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1443.000 -21.200 -1442.000 ;
    END
  END WL808
  PIN WL809
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1444.350 -21.200 -1443.350 ;
    END
  END WL809
  PIN WL810
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1446.600 -21.200 -1445.600 ;
    END
  END WL810
  PIN WL811
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1447.950 -21.200 -1446.950 ;
    END
  END WL811
  PIN WL812
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1450.200 -21.200 -1449.200 ;
    END
  END WL812
  PIN WL813
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1451.550 -21.200 -1450.550 ;
    END
  END WL813
  PIN WL814
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1453.800 -21.200 -1452.800 ;
    END
  END WL814
  PIN WL815
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1455.150 -21.200 -1454.150 ;
    END
  END WL815
  PIN WL816
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1457.400 -21.200 -1456.400 ;
    END
  END WL816
  PIN WL817
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1458.750 -21.200 -1457.750 ;
    END
  END WL817
  PIN WL818
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1461.000 -21.200 -1460.000 ;
    END
  END WL818
  PIN WL819
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1462.350 -21.200 -1461.350 ;
    END
  END WL819
  PIN WL820
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1464.600 -21.200 -1463.600 ;
    END
  END WL820
  PIN WL821
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1465.950 -21.200 -1464.950 ;
    END
  END WL821
  PIN WL822
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1468.200 -21.200 -1467.200 ;
    END
  END WL822
  PIN WL823
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1469.550 -21.200 -1468.550 ;
    END
  END WL823
  PIN WL824
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1471.800 -21.200 -1470.800 ;
    END
  END WL824
  PIN WL825
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1473.150 -21.200 -1472.150 ;
    END
  END WL825
  PIN WL826
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1475.400 -21.200 -1474.400 ;
    END
  END WL826
  PIN WL827
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1476.750 -21.200 -1475.750 ;
    END
  END WL827
  PIN WL828
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1479.000 -21.200 -1478.000 ;
    END
  END WL828
  PIN WL829
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1480.350 -21.200 -1479.350 ;
    END
  END WL829
  PIN WL830
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1482.600 -21.200 -1481.600 ;
    END
  END WL830
  PIN WL831
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1483.950 -21.200 -1482.950 ;
    END
  END WL831
  PIN WL832
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1486.200 -21.200 -1485.200 ;
    END
  END WL832
  PIN WL833
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1487.550 -21.200 -1486.550 ;
    END
  END WL833
  PIN WL834
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1489.800 -21.200 -1488.800 ;
    END
  END WL834
  PIN WL835
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1491.150 -21.200 -1490.150 ;
    END
  END WL835
  PIN WL836
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1493.400 -21.200 -1492.400 ;
    END
  END WL836
  PIN WL837
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1494.750 -21.200 -1493.750 ;
    END
  END WL837
  PIN WL838
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1497.000 -21.200 -1496.000 ;
    END
  END WL838
  PIN WL839
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1498.350 -21.200 -1497.350 ;
    END
  END WL839
  PIN WL840
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1500.600 -21.200 -1499.600 ;
    END
  END WL840
  PIN WL841
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1501.950 -21.200 -1500.950 ;
    END
  END WL841
  PIN WL842
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1504.200 -21.200 -1503.200 ;
    END
  END WL842
  PIN WL843
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1505.550 -21.200 -1504.550 ;
    END
  END WL843
  PIN WL844
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1507.800 -21.200 -1506.800 ;
    END
  END WL844
  PIN WL845
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1509.150 -21.200 -1508.150 ;
    END
  END WL845
  PIN WL846
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1511.400 -21.200 -1510.400 ;
    END
  END WL846
  PIN WL847
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1512.750 -21.200 -1511.750 ;
    END
  END WL847
  PIN WL848
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1515.000 -21.200 -1514.000 ;
    END
  END WL848
  PIN WL849
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1516.350 -21.200 -1515.350 ;
    END
  END WL849
  PIN WL850
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1518.600 -21.200 -1517.600 ;
    END
  END WL850
  PIN WL851
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1519.950 -21.200 -1518.950 ;
    END
  END WL851
  PIN WL852
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1522.200 -21.200 -1521.200 ;
    END
  END WL852
  PIN WL853
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1523.550 -21.200 -1522.550 ;
    END
  END WL853
  PIN WL854
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1525.800 -21.200 -1524.800 ;
    END
  END WL854
  PIN WL855
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1527.150 -21.200 -1526.150 ;
    END
  END WL855
  PIN WL856
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1529.400 -21.200 -1528.400 ;
    END
  END WL856
  PIN WL857
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1530.750 -21.200 -1529.750 ;
    END
  END WL857
  PIN WL858
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1533.000 -21.200 -1532.000 ;
    END
  END WL858
  PIN WL859
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1534.350 -21.200 -1533.350 ;
    END
  END WL859
  PIN WL860
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1536.600 -21.200 -1535.600 ;
    END
  END WL860
  PIN WL861
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1537.950 -21.200 -1536.950 ;
    END
  END WL861
  PIN WL862
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1540.200 -21.200 -1539.200 ;
    END
  END WL862
  PIN WL863
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1541.550 -21.200 -1540.550 ;
    END
  END WL863
  PIN WL864
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1543.800 -21.200 -1542.800 ;
    END
  END WL864
  PIN WL865
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1545.150 -21.200 -1544.150 ;
    END
  END WL865
  PIN WL866
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1547.400 -21.200 -1546.400 ;
    END
  END WL866
  PIN WL867
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1548.750 -21.200 -1547.750 ;
    END
  END WL867
  PIN WL868
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1551.000 -21.200 -1550.000 ;
    END
  END WL868
  PIN WL869
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1552.350 -21.200 -1551.350 ;
    END
  END WL869
  PIN WL870
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1554.600 -21.200 -1553.600 ;
    END
  END WL870
  PIN WL871
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1555.950 -21.200 -1554.950 ;
    END
  END WL871
  PIN WL872
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1558.200 -21.200 -1557.200 ;
    END
  END WL872
  PIN WL873
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1559.550 -21.200 -1558.550 ;
    END
  END WL873
  PIN WL874
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1561.800 -21.200 -1560.800 ;
    END
  END WL874
  PIN WL875
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1563.150 -21.200 -1562.150 ;
    END
  END WL875
  PIN WL876
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1565.400 -21.200 -1564.400 ;
    END
  END WL876
  PIN WL877
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1566.750 -21.200 -1565.750 ;
    END
  END WL877
  PIN WL878
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1569.000 -21.200 -1568.000 ;
    END
  END WL878
  PIN WL879
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1570.350 -21.200 -1569.350 ;
    END
  END WL879
  PIN WL880
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1572.600 -21.200 -1571.600 ;
    END
  END WL880
  PIN WL881
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1573.950 -21.200 -1572.950 ;
    END
  END WL881
  PIN WL882
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1576.200 -21.200 -1575.200 ;
    END
  END WL882
  PIN WL883
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1577.550 -21.200 -1576.550 ;
    END
  END WL883
  PIN WL884
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1580.350 -21.200 -1579.350 ;
    END
  END WL884
  PIN WL885
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1581.700 -21.200 -1580.700 ;
    END
  END WL885
  PIN WL886
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1583.950 -21.200 -1582.950 ;
    END
  END WL886
  PIN WL887
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1585.300 -21.200 -1584.300 ;
    END
  END WL887
  PIN WL888
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1587.550 -21.200 -1586.550 ;
    END
  END WL888
  PIN WL889
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1588.900 -21.200 -1587.900 ;
    END
  END WL889
  PIN WL890
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1591.150 -21.200 -1590.150 ;
    END
  END WL890
  PIN WL891
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1592.500 -21.200 -1591.500 ;
    END
  END WL891
  PIN WL892
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1594.750 -21.200 -1593.750 ;
    END
  END WL892
  PIN WL893
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1596.100 -21.200 -1595.100 ;
    END
  END WL893
  PIN WL894
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1598.350 -21.200 -1597.350 ;
    END
  END WL894
  PIN WL895
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1599.700 -21.200 -1598.700 ;
    END
  END WL895
  PIN WL896
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1601.950 -21.200 -1600.950 ;
    END
  END WL896
  PIN WL897
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1603.300 -21.200 -1602.300 ;
    END
  END WL897
  PIN WL898
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1605.550 -21.200 -1604.550 ;
    END
  END WL898
  PIN WL899
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1606.900 -21.200 -1605.900 ;
    END
  END WL899
  PIN WL900
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1609.150 -21.200 -1608.150 ;
    END
  END WL900
  PIN WL901
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1610.500 -21.200 -1609.500 ;
    END
  END WL901
  PIN WL902
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1612.750 -21.200 -1611.750 ;
    END
  END WL902
  PIN WL903
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1614.100 -21.200 -1613.100 ;
    END
  END WL903
  PIN WL904
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1616.350 -21.200 -1615.350 ;
    END
  END WL904
  PIN WL905
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1617.700 -21.200 -1616.700 ;
    END
  END WL905
  PIN WL906
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1619.950 -21.200 -1618.950 ;
    END
  END WL906
  PIN WL907
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1621.300 -21.200 -1620.300 ;
    END
  END WL907
  PIN WL908
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1623.550 -21.200 -1622.550 ;
    END
  END WL908
  PIN WL909
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1624.900 -21.200 -1623.900 ;
    END
  END WL909
  PIN WL910
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1627.150 -21.200 -1626.150 ;
    END
  END WL910
  PIN WL911
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1628.500 -21.200 -1627.500 ;
    END
  END WL911
  PIN WL912
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1630.750 -21.200 -1629.750 ;
    END
  END WL912
  PIN WL913
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1632.100 -21.200 -1631.100 ;
    END
  END WL913
  PIN WL914
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1634.350 -21.200 -1633.350 ;
    END
  END WL914
  PIN WL915
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1635.700 -21.200 -1634.700 ;
    END
  END WL915
  PIN WL916
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1637.950 -21.200 -1636.950 ;
    END
  END WL916
  PIN WL917
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1639.300 -21.200 -1638.300 ;
    END
  END WL917
  PIN WL918
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1641.550 -21.200 -1640.550 ;
    END
  END WL918
  PIN WL919
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1642.900 -21.200 -1641.900 ;
    END
  END WL919
  PIN WL920
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1645.150 -21.200 -1644.150 ;
    END
  END WL920
  PIN WL921
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1646.500 -21.200 -1645.500 ;
    END
  END WL921
  PIN WL922
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1648.750 -21.200 -1647.750 ;
    END
  END WL922
  PIN WL923
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1650.100 -21.200 -1649.100 ;
    END
  END WL923
  PIN WL924
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1652.350 -21.200 -1651.350 ;
    END
  END WL924
  PIN WL925
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1653.700 -21.200 -1652.700 ;
    END
  END WL925
  PIN WL926
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1655.950 -21.200 -1654.950 ;
    END
  END WL926
  PIN WL927
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1657.300 -21.200 -1656.300 ;
    END
  END WL927
  PIN WL928
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1659.550 -21.200 -1658.550 ;
    END
  END WL928
  PIN WL929
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1660.900 -21.200 -1659.900 ;
    END
  END WL929
  PIN WL930
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1663.150 -21.200 -1662.150 ;
    END
  END WL930
  PIN WL931
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1664.500 -21.200 -1663.500 ;
    END
  END WL931
  PIN WL932
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1666.750 -21.200 -1665.750 ;
    END
  END WL932
  PIN WL933
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1668.100 -21.200 -1667.100 ;
    END
  END WL933
  PIN WL934
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1670.350 -21.200 -1669.350 ;
    END
  END WL934
  PIN WL935
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1671.700 -21.200 -1670.700 ;
    END
  END WL935
  PIN WL936
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1673.950 -21.200 -1672.950 ;
    END
  END WL936
  PIN WL937
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1675.300 -21.200 -1674.300 ;
    END
  END WL937
  PIN WL938
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1677.550 -21.200 -1676.550 ;
    END
  END WL938
  PIN WL939
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1678.900 -21.200 -1677.900 ;
    END
  END WL939
  PIN WL940
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1681.150 -21.200 -1680.150 ;
    END
  END WL940
  PIN WL941
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1682.500 -21.200 -1681.500 ;
    END
  END WL941
  PIN WL942
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1684.750 -21.200 -1683.750 ;
    END
  END WL942
  PIN WL943
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1686.100 -21.200 -1685.100 ;
    END
  END WL943
  PIN WL944
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1688.350 -21.200 -1687.350 ;
    END
  END WL944
  PIN WL945
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1689.700 -21.200 -1688.700 ;
    END
  END WL945
  PIN WL946
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1691.950 -21.200 -1690.950 ;
    END
  END WL946
  PIN WL947
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1693.300 -21.200 -1692.300 ;
    END
  END WL947
  PIN WL948
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1695.550 -21.200 -1694.550 ;
    END
  END WL948
  PIN WL949
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1696.900 -21.200 -1695.900 ;
    END
  END WL949
  PIN WL950
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1699.150 -21.200 -1698.150 ;
    END
  END WL950
  PIN WL951
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1700.500 -21.200 -1699.500 ;
    END
  END WL951
  PIN WL952
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1702.750 -21.200 -1701.750 ;
    END
  END WL952
  PIN WL953
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1704.100 -21.200 -1703.100 ;
    END
  END WL953
  PIN WL954
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1706.350 -21.200 -1705.350 ;
    END
  END WL954
  PIN WL955
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1707.700 -21.200 -1706.700 ;
    END
  END WL955
  PIN WL956
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1709.950 -21.200 -1708.950 ;
    END
  END WL956
  PIN WL957
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1711.300 -21.200 -1710.300 ;
    END
  END WL957
  PIN WL958
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1713.550 -21.200 -1712.550 ;
    END
  END WL958
  PIN WL959
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1714.900 -21.200 -1713.900 ;
    END
  END WL959
  PIN WL960
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1717.150 -21.200 -1716.150 ;
    END
  END WL960
  PIN WL961
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1718.500 -21.200 -1717.500 ;
    END
  END WL961
  PIN WL962
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1720.750 -21.200 -1719.750 ;
    END
  END WL962
  PIN WL963
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1722.100 -21.200 -1721.100 ;
    END
  END WL963
  PIN WL964
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1724.350 -21.200 -1723.350 ;
    END
  END WL964
  PIN WL965
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1725.700 -21.200 -1724.700 ;
    END
  END WL965
  PIN WL966
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1727.950 -21.200 -1726.950 ;
    END
  END WL966
  PIN WL967
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1729.300 -21.200 -1728.300 ;
    END
  END WL967
  PIN WL968
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1731.550 -21.200 -1730.550 ;
    END
  END WL968
  PIN WL969
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1732.900 -21.200 -1731.900 ;
    END
  END WL969
  PIN WL970
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1735.150 -21.200 -1734.150 ;
    END
  END WL970
  PIN WL971
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1736.500 -21.200 -1735.500 ;
    END
  END WL971
  PIN WL972
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1738.750 -21.200 -1737.750 ;
    END
  END WL972
  PIN WL973
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1740.100 -21.200 -1739.100 ;
    END
  END WL973
  PIN WL974
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1742.350 -21.200 -1741.350 ;
    END
  END WL974
  PIN WL975
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1743.700 -21.200 -1742.700 ;
    END
  END WL975
  PIN WL976
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1745.950 -21.200 -1744.950 ;
    END
  END WL976
  PIN WL977
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1747.300 -21.200 -1746.300 ;
    END
  END WL977
  PIN WL978
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1749.550 -21.200 -1748.550 ;
    END
  END WL978
  PIN WL979
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1750.900 -21.200 -1749.900 ;
    END
  END WL979
  PIN WL980
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1753.150 -21.200 -1752.150 ;
    END
  END WL980
  PIN WL981
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1754.500 -21.200 -1753.500 ;
    END
  END WL981
  PIN WL982
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1756.750 -21.200 -1755.750 ;
    END
  END WL982
  PIN WL983
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1758.100 -21.200 -1757.100 ;
    END
  END WL983
  PIN WL984
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1760.350 -21.200 -1759.350 ;
    END
  END WL984
  PIN WL985
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1761.700 -21.200 -1760.700 ;
    END
  END WL985
  PIN WL986
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1763.950 -21.200 -1762.950 ;
    END
  END WL986
  PIN WL987
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1765.300 -21.200 -1764.300 ;
    END
  END WL987
  PIN WL988
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1767.550 -21.200 -1766.550 ;
    END
  END WL988
  PIN WL989
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1768.900 -21.200 -1767.900 ;
    END
  END WL989
  PIN WL990
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1771.150 -21.200 -1770.150 ;
    END
  END WL990
  PIN WL991
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1772.500 -21.200 -1771.500 ;
    END
  END WL991
  PIN WL992
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1774.750 -21.200 -1773.750 ;
    END
  END WL992
  PIN WL993
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1776.100 -21.200 -1775.100 ;
    END
  END WL993
  PIN WL994
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1778.900 -21.200 -1777.900 ;
    END
  END WL994
  PIN WL995
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1780.250 -21.200 -1779.250 ;
    END
  END WL995
  PIN WL996
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1782.500 -21.200 -1781.500 ;
    END
  END WL996
  PIN WL997
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1783.850 -21.200 -1782.850 ;
    END
  END WL997
  PIN WL998
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1786.100 -21.200 -1785.100 ;
    END
  END WL998
  PIN WL999
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1787.450 -21.200 -1786.450 ;
    END
  END WL999
  PIN WL1000
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1789.700 -21.200 -1788.700 ;
    END
  END WL1000
  PIN WL1001
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1791.050 -21.200 -1790.050 ;
    END
  END WL1001
  PIN WL1002
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1793.300 -21.200 -1792.300 ;
    END
  END WL1002
  PIN WL1003
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1794.650 -21.200 -1793.650 ;
    END
  END WL1003
  PIN WL1004
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1796.900 -21.200 -1795.900 ;
    END
  END WL1004
  PIN WL1005
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1798.250 -21.200 -1797.250 ;
    END
  END WL1005
  PIN WL1006
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1800.500 -21.200 -1799.500 ;
    END
  END WL1006
  PIN WL1007
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1801.850 -21.200 -1800.850 ;
    END
  END WL1007
  PIN WL1008
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1804.100 -21.200 -1803.100 ;
    END
  END WL1008
  PIN WL1009
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1805.450 -21.200 -1804.450 ;
    END
  END WL1009
  PIN WL1010
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1807.700 -21.200 -1806.700 ;
    END
  END WL1010
  PIN WL1011
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1809.050 -21.200 -1808.050 ;
    END
  END WL1011
  PIN WL1012
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1811.300 -21.200 -1810.300 ;
    END
  END WL1012
  PIN WL1013
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1812.650 -21.200 -1811.650 ;
    END
  END WL1013
  PIN WL1014
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1814.900 -21.200 -1813.900 ;
    END
  END WL1014
  PIN WL1015
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1816.250 -21.200 -1815.250 ;
    END
  END WL1015
  PIN WL1016
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1818.500 -21.200 -1817.500 ;
    END
  END WL1016
  PIN WL1017
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1819.850 -21.200 -1818.850 ;
    END
  END WL1017
  PIN WL1018
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1822.100 -21.200 -1821.100 ;
    END
  END WL1018
  PIN WL1019
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1823.450 -21.200 -1822.450 ;
    END
  END WL1019
  PIN WL1020
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1825.700 -21.200 -1824.700 ;
    END
  END WL1020
  PIN WL1021
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1827.050 -21.200 -1826.050 ;
    END
  END WL1021
  PIN WL1022
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1829.300 -21.200 -1828.300 ;
    END
  END WL1022
  PIN WL1023
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met3 ;
        RECT -23.200 -1830.650 -21.200 -1829.650 ;
    END
  END WL1023
  PIN vssd1
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -23.200 26.000 -21.200 28.000 ;
        RECT 226.000 26.000 228.000 28.000 ;
        RECT -23.200 -1868.000 228.000 -1866.000 ;
    END
  END vssd1
  PIN vccd1
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT -21.000 31.000 -19.000 33.000 ;
        RECT -7.950 31.000 -6.950 32.500 ;
        RECT 217.800 31.000 218.800 32.500 ;
        RECT 226.000 -1873.000 228.000 33.000 ;
      LAYER via2 ;
        RECT -20.500 31.500 -19.500 32.500 ;
        RECT -7.850 31.600 -7.050 32.400 ;
        RECT 217.900 31.600 218.700 32.400 ;
        RECT 226.500 31.500 227.500 32.500 ;
        RECT 226.900 -1855.600 227.400 -1855.150 ;
        RECT 226.500 -1872.500 227.500 -1871.500 ;
      LAYER met3 ;
        RECT -23.200 31.000 228.000 33.000 ;
        RECT 226.000 -1855.750 227.500 -1855.000 ;
        RECT -23.200 -1873.000 228.000 -1871.000 ;
    END
  END vccd1
  OBS
      LAYER li1 ;
        RECT -11.270 -1864.100 218.050 22.080 ;
      LAYER met1 ;
        RECT -11.270 -1864.100 223.000 22.170 ;
      LAYER met2 ;
        RECT -21.000 -1873.000 223.000 31.000 ;
      LAYER met3 ;
        RECT -21.200 -1855.750 226.000 28.000 ;
  END
END full_sram
END LIBRARY

